package shared_pkg;
 logic test_finished;
 integer error_counter=0;
 integer Correct_counter=0;
endpackage : shared_pkg